module display_tb;
    initial begin
        $display("display tb");
    end
endmodule
