module debounce(src, dst);
    input  src;
    output dst;
endmodule
