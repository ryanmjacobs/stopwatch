module top;
	module clkdiv();
	module display();
endmodule
