module display(seconds);
    input seconds;
endmodule
