module top_tb;
    initial begin
        #1 $display("top tb");
    end
endmodule
