module debounce_tb;
    initial begin
        $display("debounce tb");
    end
endmodule
